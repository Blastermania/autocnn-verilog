// Top-level CNN module
module cnn_top (
    input wire clk, reset,
    input wire [1*16-1:0] input_data,
    output wire [10*16-1:0] output_data
);

// TODO: Instantiate conv2d, relu, maxpool, fc modules here

endmodule